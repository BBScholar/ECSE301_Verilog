

module s_adder(
	input x, y, kin, en,
	output u, kout
);

always begin

end


endmodule
