

module testbench2();

    wire rst, clk;
    wire [2:0] ls;
    wire [2:0] ls;


endmodule
